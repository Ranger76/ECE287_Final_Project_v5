library ieee;
use ieee.std_logic_1164.all;

package state_type is
	type state_type is (STATE_1, STATE_2, STATE_3, STATE_4, STATE_5, STATE_6, STATE_Collide_Check);
end package state_type;
